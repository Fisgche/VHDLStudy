LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Decodificador_74LS138 IS 
PORT(
	E: IN STD_LOGIC_VECTOR(3 DOWNTO 1);
	A: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	O: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END ENTITY;

--------------------------

ARCHITECTURE arch OF Decodificador_74LS138 IS
SIGNAL aux : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	WITH A SELECT 
		aux <= "11111110" WHEN "000",
			"11111101" WHEN "001",
			"11111011" WHEN "010",
			"11110111" WHEN "011",
			"11101111" WHEN "100",
			"11011111" WHEN "101",
			"10111111" WHEN "110",
			"01111111" WHEN "111";
	O <= aux WHEN e = "100" ELSE "00000000";
END arch;
